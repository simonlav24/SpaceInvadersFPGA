// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen FWbruary  2021  
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	ScoreBoardDigits	(	
					input	logic	clk,
					input	logic	resetN,
					input   logic	[10:0] offsetX,// offset from top left  position 
					input   logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
                    
                    input logic [3:0] digit0,
                    input logic [3:0] digit1,
                    input logic [3:0] digit2,
                    input logic [3:0] digit3,
                    input logic [3:0] digit4,
					
					output logic	drawingRequest, //output that the pixel should be dispalyed 
					output logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hde ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */

//logic [10:0] monster_shootX_ins;
//logic [10:0] monster_shootY_ins;

//int counterX = 3;
//int counterY = 0; 

//logic [1:0] monster_type = 2'b00;

// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 

//
//logic [0:4] [0:9] MazeBiMapMask;
//
//logic [0:4] [0:4] MazeInit = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000};

//////num////Y//////X
bit [0:15] [0:15] [0:15] object_colors  = {
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0001100001111000,
16'b 0001100001111000,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0001111000011000,
16'b 0001111000011000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000000000,
16'b 0000000000000000},


																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0001111110000000,
16'b 0001111110000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0111111111111000,
16'b 0111111111111000,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0000000001111110,
16'b 0000000001111110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111111000000000,
16'b 0111111000000000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0001111111111110,
16'b 0001111111111110,
16'b 0000000001111000,
16'b 0000000001111000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000011110,
16'b 0000000000011110,
16'b 0110000000011110,
16'b 0110000000011110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000000111111000,
16'b 0000000111111000,
16'b 0000011111111000,
16'b 0000011111111000,
16'b 0001111001111000,
16'b 0001111001111000,
16'b 0111100001111000,
16'b 0111100001111000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0000000001111000,
16'b 0000000001111000,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0111111111111000,
16'b 0111111111111000,
16'b 0110000000000000,
16'b 0110000000000000,
16'b 0111111111111000,
16'b 0111111111111000,
16'b 0000000000011110,
16'b 0000000000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111100000000000,
16'b 0111100000000000,
16'b 0111111111111000,
16'b 0111111111111000,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0000000001111000,
16'b 0000000001111000,
16'b 0000000111100000,
16'b 0000000111100000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0000011110000000,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000000000000000,
16'b 0000000000000000},
																	
{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0111100000011110,
16'b 0001111111111110,
16'b 0001111111111110,
16'b 0000000000011110,
16'b 0000000000011110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000000000000000,
16'b 0000000000000000},

{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000000000,
16'b 0000000000000000},


{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000000000,
16'b 0000000000000000},

{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000000000,
16'b 0000000000000000},


{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000000000,
16'b 0000000000000000},

{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000000000,
16'b 0000000000000000},

{16'b 0000000000000000,
16'b 0000000000000000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0111111111111110,
16'b 0001111111111000,
16'b 0001111111111000,
16'b 0000011111100000,
16'b 0000011111100000,
16'b 0000000000000000,
16'b 0000000000000000}
} ; 

logic [7:0] digit_color = 8'hff ; //set the color of the digit 

logic [3:0] num_type;
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		//MazeBiMapMask <= MazeInit;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if (InsideRectangle == 1'b1 ) begin 
			if (offsetX[8:4] == 		5'b00000)
				num_type <= digit4;
			else if(offsetX[8:4] == 5'b00001)
				num_type <= digit3;
			else if(offsetX[8:4] == 5'b00010)
				num_type <= digit2;
			else if(offsetX[8:4] == 5'b00011)
				num_type <= digit1;
			else if(offsetX[8:4] == 5'b00100)
				num_type <= digit0;
         if(object_colors[num_type][offsetY[3:0]][offsetX[3:0]] == 1) begin
             RGBout <= digit_color;
         end
		end
	end
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap  
endmodule

