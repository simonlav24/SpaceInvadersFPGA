// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen FWbruary  2021  
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	HartsMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket \
					input logic collision_missile,
					input logic [10:0] missileX,
					input logic [10:0] missileY,
					
					input logic [10:0] topleftX,
					input logic [10:0] topleftY,
					input logic startOfFrame,

					output logic [10:0] monster_shootX,
					output logic [10:0] monster_shootY,
					
					output logic	drawingRequest, //output that the pixel should be dispalyed 
					output logic	[7:0] RGBout,  //rgb value from the bitmap 
					
					output logic win
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hde ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */

logic [10:0] monster_shootX_ins;
logic [10:0] monster_shootY_ins;

int counterX = 3;
int counterY = 0; 

int anim_counter = 0;
logic anim_type = 1'b0;

logic [2:0] monster_type = 3'b000;

// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 

int alienCounter = 0;

logic [0:4] [0:9]  MazeBiMapMask;

logic [0:4] [0:9] MazeInit = 
{10'b	1111111111,
10'b	1111111111,
10'b	1111111111,
10'b	1111111111,
10'b	1111111111};

 
 logic [0:7] [0:31] [0:31] [7:0]  object_colors  = {
 // alien 1A
{  {8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}
},

{// alien 1B
   {8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'h1f,8'h1f,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}
},
// alien 2A
{  {8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}
},

{// alien 2B
   {8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hea,8'hea,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hea,8'hea,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}
},
{	// alien 3A
   {8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}
},

{  //alien 3B
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'he4,8'he4,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}

},

{ // alien 4A
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}

},

{/// alien 4B
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hef,8'hef,8'hef,8'hef,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde},
	{8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde,8'hde}
}
};
 
logic noMoreAliens = 1'b0;
 
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBiMapMask <= MazeInit;
		counterX <= 0;
		counterY <= 0;
		monster_type <= 3'b00;
		anim_counter <= 0;
		noMoreAliens <= 1'b0;
		alienCounter <= 0;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if (InsideRectangle == 1'b1 ) begin 
		   if (MazeBiMapMask[offsetY[8:5] ][offsetX[8:5]] == 1'b1 ) begin// if in 32 grid
				
				if 	 (offsetY[8:5] == 2'b00)
					monster_type <= 3'b000 | anim_type;
				else if(offsetY[8:5] == 2'b01)
					monster_type <= 3'b000 | anim_type;
				else if(offsetY[8:5] == 2'b10)
					monster_type <= 3'b110 | anim_type;
				else if(offsetY[8:5] == 2'b11)
					monster_type <= 3'b100 | anim_type;
				else if(offsetY[8:5] == 3'b100)
					monster_type <= 3'b010 | anim_type;
					
				RGBout <= object_colors[monster_type][offsetY[4:0]][offsetX[4:0]] ;
			end
		end
		
		if (collision_missile == 1'b1) begin
			MazeBiMapMask[offsetY[8:5]] [offsetX[8:5]] = 1'b0;
			alienCounter <= alienCounter + 1;
		end
		
		if (alienCounter >= 50)
			noMoreAliens <= 1'b1;
		
		if (startOfFrame == 1'b1) begin
		
			anim_counter <= anim_counter + 1;
			if(anim_counter == 30) begin
				anim_counter <= 0;
				anim_type <= ~anim_type;
			end
		
			counterX <= counterX + 1;
			if (counterX > 9) begin
				counterX <= 0;
				counterY <= counterY + 1;
				if (counterY > 4)
					counterY <= 0;
			end
				
		
			if (MazeBiMapMask[counterY][counterX] == 1'b1) begin
				// get monster position
				monster_shootX_ins <= topleftX + 16 + 32 * counterX;
				monster_shootY_ins <= topleftY + 16 + 32 * counterY;
				
			end
		end
		
	
		
		
	end
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap  
assign monster_shootX = monster_shootX_ins;
assign monster_shootY = monster_shootY_ins;
assign win = noMoreAliens;
endmodule

