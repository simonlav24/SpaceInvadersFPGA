// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen FWbruary  2021  
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	end_screen	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket \
					
					input logic [10:0] topleftX,
					input logic [10:0] topleftY,
					input logic startOfFrame,
					
					input logic win,
					
					output logic	drawingRequest, //output that the pixel should be dispalyed 
					output logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hde ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 
int counter= 0;

logic [0:1] [0:5] [0:64]  title =
{
{
65'b  01111100011100001110110000111100000001111000100010001111000100111,
65'b  10000100000010001001001001000010000010000100100010010000100101000,
65'b  10000100011110001001001001111110000010000100100010011111100110000,
65'b  01111100100010001001001001000000000010000100010100010000000100000,
65'b  00000100011111001001001000111110000001111000001000001111100100000,
65'b  11111000000000000000000000000000000000000000000000000000000000000
},
{
65'b  00000000001000100011110001000100000100000100100111100010000000000,
65'b  00000000001000100100001001000100000100100100100100010010000000000,
65'b  00000000001000100100001001000100000100100100100100010010000000000,
65'b  00000000000111100100001001000100000101010100100100010010000000000,
65'b  00000000000000100011110000111100000010001000100100010000000000000,
65'b  00000000001111000000000000000000000000000000000000000010000000000
}
};

 
//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if (InsideRectangle == 1'b1 ) begin 
		   if (title[win][offsetY[10:2] ][offsetX[10:2]] == 1'b1 ) begin// if in 32 grid
				
				
				RGBout <= 8'hff;
			end
		end
		
		if (startOfFrame == 1'b1) begin
			counter = counter + 1;
		end

	end
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap  
endmodule

